parameter C = 5'b00001;
parameter Csharp = 5'b00010;
parameter D = 5'b00011;
parameter Dsharp = 5'b00100;
parameter E = 5'b00101;
parameter F = 5'b00110;
parameter Fsharp = 5'b00111;
parameter G = 5'b01000;
parameter Gsharp = 5'b01001;
parameter A = 5'b01010;
parameter Asharp = 5'b01011;
parameter B = 5'01100;
parameter C2 = 5'01101;
parameter Csharp2 = 5'01110;
parameter D2 = 5'01111;
parameter Dsharp2 = 5'b10000;
parameter E2 = 5'b10001;
parameter F2 = 5'b10010;
parameter Fsharp2 = 5'b10011;
parameter G2 = 5'b10100;
parameter Gsharp2 = 5'b10101;
parameter A2 = 5'b10110;
parameter Asharp2 = 5'b10111;
parameter B2 = 5'b11000;
parameter C3 = 5'b11001;

parameter tSINE = 3'b000, tSQUARE = 3'b001, tSAW = 3'b010;

parameter hexA = 6'd1;
parameter hexB = 6'd2;
parameter hexC = 6'd3;
parameter hexD = 6'd4;
parameter hexE = 6'd5;
parameter hexF = 6'd6;
parameter hexG = 6'd7;
parameter hexH = 6'd8;
parameter hexI = 6'd9;
parameter hexJ = 6'd10;
parameter hexK = 6'd11;
parameter hexL = 6'd12;
parameter hexM = 6'd13;
parameter hexN = 6'd14;
parameter hexO = 6'd15;
parameter hexP = 6'd16;
parameter hexQ = 6'd17;
parameter hexR = 6'd18;
parameter hexS = 6'd19;
parameter hexT = 6'd20;
parameter hexU = 6'd21;
parameter hexV = 6'd22;
parameter hexW = 6'd23;
parameter hexX = 6'd24;
parameter hexY = 6'd25;
parameter hexZ = 6'd26;

parameter hex0 = 6'd27;
parameter hex1 = 6'd28;
parameter hex2 = 6'd29;
parameter hex3 = 6'd30;
parameter hex4 = 6'd31;
parameter hex5 = 6'd32;
parameter hex6 = 6'd33;
parameter hex7 = 6'd34;
parameter hex8 = 6'd35;
parameter hex9 = 6'd36;