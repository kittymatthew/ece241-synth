parameter C = 5'b00001;
parameter Csharp = 5'b00010;
parameter D = 5'b00011;
parameter Dsharp = 5'b00100;
parameter E = 5'b00101;
parameter F = 5'b00110;
parameter Fsharp = 5'b00111;
parameter G = 5'b01000;
parameter Gsharp = 5'b01001;
parameter A = 5'b01010;
parameter Asharp = 5'b01011;
parameter B = 5'01100;
parameter C2 = 5'01101;
parameter Csharp2 = 5'01110;
parameter D2 = 5'01111;
parameter Dsharp2 = 5'b10000;
parameter E2 = 5'b10001;
parameter F2 = 5'b10010;
parameter Fsharp2 = 5'b10011;
parameter G2 = 5'b10100;
parameter Gsharp2 = 5'b10101;
parameter A2 = 5'b10110;
parameter Asharp2 = 5'b10111;
parameter B2 = 5'b11000;
parameter C3 = 5'b11001;

parameter tSINE = 3'b000, tSQUARE = 3'b001, tSAW = 3'b010;