module waveform_gen (TYPE, NOTE, OUT, clock, enable, reset);
    input [2:0] TYPE;
    input [4:0] NOTE;
    input clock, enable, reset;

    wire [31:0] SINE, SQUARE, SAW;
    reg [31:0] BUFFER;
    output reg [31:0] OUT;

    sine_gen sine_generator (NOTE, SINE, clock, reset);
    square_gen square_gen (NOTE, SQUARE, clock, reset);
    saw_gen saw_gen (NOTE, SAW, clock, reset);

    parameter tSINE = 3'b000, tSQUARE = 3'b001, tSAW = 3'b010;

    always @ (*) begin
        case (TYPE) // Output the approriate waveform type
            tSINE: begin BUFFER = SINE; end
            tSQUARE: begin BUFFER = SQUARE; end
            tSAW: begin BUFFER = SAW; end
            default: begin BUFFER = 32'b0; end
        endcase
    end

    always @ (posedge clock, posedge reset) begin
        if (reset) begin // Reset on reset signal
            OUT <= 32'b0; 
        end
        else if (enable) begin OUT <= BUFFER; end // Only output when enable is high
        else begin OUT <= OUT; end
    end
endmodule

module sine_gen (NOTE, OUT, clock, reset);
    input [4:0] NOTE; // 5-bit number representing which note frequency we should generate 
    input clock, reset; // Clock and reset signals

    output reg [31:0] OUT; // 32-bit unsigned output
    reg [31:0] COUNT, STEP; // Counter and step values, see note below

    reg [31:0] SINE_LUT [0:1023]; // 1024-value 32-bit sine lookup table - so we don't have to calculate sine ourselves

    /* 
        To save 1024 lines of code, we directly read sine_lookup.hex into the SINE_LUT registers. 
        Each line of sine_lookup.hex is a hexadecimal value between 0 and 2^32-1, mapped to the shape of a sine wave.
        The values were generated by https://www.daycounter.com/Calculators/Sine-Generator-Calculator.phtml.
    */
    initial begin
        $readmemh("sine_lookup.hex", SINE_LUT, 0, 1023);
    end

    // The waveform can generate two full octaves, see note below
    parameter C = 5'b00001;
    parameter Csharp = 5'b00010;
    parameter D = 5'b00011;
    parameter Dsharp = 5'b00100;
    parameter E = 5'b00101;
    parameter F = 5'b00110;
    parameter Fsharp = 5'b00111;
    parameter G = 5'b01000;
    parameter Gsharp = 5'b01001;
    parameter A = 5'b01010;
    parameter Asharp = 5'b01011;
    parameter B = 5'b01100;
    parameter C2 = 5'b01101;
    parameter Csharp2 = 5'b01110;
    parameter D2 = 5'b01111;
    parameter Dsharp2 = 5'b10000;
    parameter E2 = 5'b10001;
    parameter F2 = 5'b10010;
    parameter Fsharp2 = 5'b10011;
    parameter G2 = 5'b10100;
    parameter Gsharp2 = 5'b10101;
    parameter A2 = 5'b10110;
    parameter Asharp2 = 5'b10111;
    parameter B2 = 5'b11000;
    parameter C3 = 5'b11001;

    /* 
        The frequency we output is determined based on how 'fast' we traverse through the sine wave.
        We change the speed we traverse through the sine wave based on how many entries of the lookup table we travel through.
        We can calculate this using: increment = (f_out * 2^32) / f_clk
        However, because we want to synthesize this code, we try to avoid using division, so we hard-coded the step values for two full octaves.
        We round the step to the nearest whole number, but because they are so large, this is not noticeable
    */
    always @ (*) begin
        case (NOTE)
            C:       STEP = 32'd22474; // 261.63 Hz
            Csharp:  STEP = 32'd23809; // 277.18 Hz
            D:       STEP = 32'd25225; // 293.66 Hz
            Dsharp:  STEP = 32'd26726; // 311.13 Hz
            E:       STEP = 32'd28315; // 329.63 Hz
            F:       STEP = 32'd29999; // 349.23 Hz
            Fsharp:  STEP = 32'd31782; // 369.99 Hz
            G:       STEP = 32'd33673; // 392.00 Hz
            Gsharp:  STEP = 32'd35674; // 415.30 Hz
            A:       STEP = 32'd37796; // 440.00 Hz
            Asharp:  STEP = 32'd40043; // 466.16 Hz
            B:       STEP = 32'd42424; // 493.88 Hz
            C2:      STEP = 32'd44947; // 523.25 Hz
            Csharp2: STEP = 32'd47620; // 554.37 Hz
            D2:      STEP = 32'd50451; // 587.33 Hz
            Dsharp2: STEP = 32'd53451; // 622.25 Hz
            E2:      STEP = 32'd56630; // 659.26 Hz
            F2:      STEP = 32'd59997; // 698.46 Hz
            Fsharp2: STEP = 32'd63565; // 739.99 Hz
            G2:      STEP = 32'd67344; // 783.99 Hz
            Gsharp2: STEP = 32'd71349; // 830.61 Hz
            A2:      STEP = 32'd75591; // 880.00 Hz
            Asharp2: STEP = 32'd80087; // 932.33 Hz
            B2:      STEP = 32'd84849; // 987.77 Hz
            C3:      STEP = 32'd89901; // 1046.59 Hz
            default: STEP = 32'd0;
        endcase
    end

    // The generation is based off of a phase-accumulator: see https://www.analog.com/en/resources/analog-dialogue/articles/all-about-direct-digital-synthesis.html.

    wire [31:0] next_count = COUNT + STEP; // next_count is the next count we need to progress to
    wire [9:0] next_address = next_count[31:22]; // Only use the upper bits of next_count - this saves us from having to use a sine LUT with tens of thousands of entries

    always @ (posedge clock, posedge reset) begin
        if (reset) begin // Reset the signals on reset
            COUNT <= 32'b0; 
            OUT <= 32'b0; 
        end else begin
            COUNT <= next_count; // Increment the count by next_count, which determines the frequency we are playing
            OUT <= SINE_LUT[next_address]; // Output the appropriate sine value
        end
    end
endmodule

// Square wave generator - will be implemented later, time permitting
module square_gen (FREQUENCY, OUT, clock, reset);
    input [4:0] FREQUENCY;
    input clock, reset;

    output [31:0] OUT;
endmodule

// Sawtooth wave generator - will be implmented later, time permitting
module saw_gen (FREQUENCY, OUT, clock, reset);
    input [4:0] FREQUENCY;
    input clock, reset;

    output [31:0] OUT;
endmodule